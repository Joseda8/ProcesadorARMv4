module Negative #(parameter N = 3)(input logic r, output logic z);

	assign z = r;

endmodule
